`default_nettype none
`define default_netname none

// User IN
`define UI_IN_CLOCK         0
`define UI_IN_RESET         1
`define UI_IN_SCI_CSN       2
`define UI_IN_SCI_REQ       3
`define UI_IN_LOAD_IN       4
`define UI_IN_LOAD_VALUE_IN 5
`define UI_IN_SHIFT_OUT     6
`define UI_IN_START         7

// User OUT
`define UO_OUT_SCI_RESP         0
`define UO_OUT_SCI_ACK          1
`define UO_OUT_SHIFT_VALUE_OUT  2
`define UO_OUT_READY            3
`define UO_OUT_DONE             4

module tt_um_scorbetta_goa
(
    input wire [7:0]    ui_in, // Dedicated inputs
    output wire [7:0]   uo_out, // Dedicated outputs
    input wire [7:0]    uio_in, // IOs: Input path
    output wire [7:0]   uio_out, // IOs: Output path
    output wire [7:0]   uio_oe, // IOs: Enable path (active high: 0=input, 1=output)
    input wire          ena, // will go high when the design is enabled
    input wire          clk, // clock
    input wire          rst_n // reset_n - low to reset
);

    wire [7:0]  counter;
    wire        tt_rstn_i;
    wire        fpga_rstn_i;

    // Keep the design under reset if not enabled
    assign tt_rstn_i    = ena & rst_n;
    assign fpga_rstn_i  = ena & ui_in[`UI_IN_RESET];

    // Use main clock to check power
    COUNTER #(
        .WIDTH  (8)
    )
    COUNTER (
        .CLK        (clk),
        .RSTN       (tt_rstn_i),
        .EN         (ena),
        .VALUE      (counter),
        .OVERFLOW   () // Unused
    );

    // Check three MSBs
    assign uo_out[7:5] = counter[7:5];

    // User design uses a custom clock, generated by remote FPGA
    NEURON_WRAPPER NEURON_WRAPPER (
        .CLK                (ui_in[`UI_IN_CLOCK]),
        .RSTN               (fpga_rstn_i),
        .SCI_CSN            (ui_in[`UI_IN_SCI_CSN]),
        .SCI_REQ            (ui_in[`UI_IN_SCI_REQ]),
        .SCI_RESP           (uo_out[`UO_OUT_SCI_RESP]),
        .SCI_ACK            (uo_out[`UO_OUT_SCI_ACK]),
        .LOAD_IN            (ui_in[`UI_IN_LOAD_IN]),
        .LOAD_VALUE_IN      (ui_in[`UI_IN_LOAD_VALUE_IN]),
        .SHIFT_OUT          (ui_in[`UI_IN_SHIFT_OUT]),
        .SHIFT_VALUE_OUT    (uo_out[`UO_OUT_SHIFT_VALUE_OUT]),
        .READY              (uo_out[`UO_OUT_READY]),
        .START              (ui_in[`UI_IN_START]),
        .DONE               (uo_out[`UO_OUT_DONE])
    );

    // Bidirectional pins are not used
    assign uio_out  = 0;
    assign uio_oe   = 0;
endmodule

`default_nettype wire
